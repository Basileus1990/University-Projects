2023-01-15_22:36:52
 �������������������������������   6�&1�@        �           ����      $�       ���"  h  ����      �?    ���� ���������������������������������̎  �   ����           ���� ������������������������������� ������������������������������� ������������������������������� ����������������������������������a  L   ����           ����2023-01-15_22:42:02
 �������������������������������   �23333 @        K  �  2   ����      $�       ���  h  ����      �?    �������(  �   ����           ������̹  ;  ����           ���� ����������������������������������@  �   ����           �������H  u  ����           �������=  2   ����           ������̒  �  ����           ����2023-01-15_22:42:18
 �������������������������������   ���� 0'@        D  �  2   ����      $�       ���[  h  ����      �?    ��������   W  ����           �������!  F   ����           ���� ������������������������������� �����������������������������������   �  ����           ��������   �   ����           ���� �������������������������������2023-01-15_22:43:14
 �������������������������������   �23333$@ޭG�z@�          ����      $�       ���^  h  ����      �?    ���� ������������������������������� ������������������������������� ������������������������������� ���������������������������������̂  �  ����           �������y  �   ����           ������̖  H  ����           ����2023-01-15_22:45:19
 �������������������������������   C��K�@�+�Y@L           ����      $�       ���@  h  ����      �?    ���� ������������������������������� ������������������������������� ������������������������������� ������������������������������� ������������������������������� ������������������������������� �������������������������������2023-01-15_22:48:46
 �������������������������������   �W9��v"@        N  N      ���̌z�Ga@       ����   h  ����      �?    �������<     ����           ���� ������������������������������� ������������������������������� ����������������������������������p  m  ����           �������=  �   ����           ���� �������������������������������2023-01-15_22:52:15
 �������������������������������   ��Zd�@          �  d   ����      $�       ����   h  �����(\���@    �������_  F   �����(\���@   �������F  �  �������Q��?   ���� ����������������������������������`  �   �����(\���@   ���� ����������������������������������:    �������Q��?   �������  l  �������Q��?   ����2023-01-15_22:52:26
 �������������������������������   ���Q�2@        2  2  �   ����B�~j��.@       ���  h  ����_���(\@    ���� ���������������������������������̾   q  �������Q��?   �������  �   ���̾��Q��?   �������  !  ���̾��Q��?   ���� ����������������������������������6     ���̾��Q��?   ��������   g  �������Q��?   ����2023-01-15_22:52:42
 �������������������������������   {�&1��?        &           ����      $�       ���@  h  ����      �?    ���� ������������������������������� ������������������������������� ������������������������������� ������������������������������� ������������������������������� ������������������������������� �������������������������������